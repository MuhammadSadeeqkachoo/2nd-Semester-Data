* D:\2nd semester\CIRCUIT AND SYSTEMS 1 LAB\lab 12\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Jul 02 17:26:31 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
